* C:\Users\saisr\eSim-Workspace\esim_1\esim_1.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 5/14/2021 3:12:28 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U4  in1 in2 Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_2		
v1  in1 GND pulse		
R1  out1 GND resistor		
U3  in1 plot_v1		
R2  out2 GND resistor		
R3  out3 GND resistor		
R4  out4 GND resistor		
v2  in2 GND pulse		
U2  in2 plot_v1		
U10  out1 plot_v1		
U7  out2 plot_v1		
U11  out3 plot_v1		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ lfsr		
U5  Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ out1 out2 out3 out4 dac_bridge_4		

.end
